/*
    Unsigned 8 bit multipler with testbench
*/

module testbench(
);
    reg clk; 

    always
    begin
        clk <= 1; # 5; clk <= 0; # 5;
    end 

    wire [63:0] nxtProduct;
    reg  [63:0]  Product;
    reg  [32:0]   op1; 
    reg  [32:0]   op2; 
    wire [63:0] nxtChkProduct;
    reg  [63:0] chkProduct; 
    reg fail; 

    initial begin
        op1 <= 0;
        op2 <= 0;
        Product <= 0;
        chkProduct <= 0;
        clk <= 0; 
        fail <=0;
    end 

    always @(posedge clk) begin 
        Product <= nxtProduct;
        op1 <= op1 +1; 
        if(op1 === 256) begin
            op2 <= op2+1;
            op1 <= 0; 
        end
        chkProduct <= nxtChkProduct; 
     end

    multipler mul(op1[31:0],op2[31:0],nxtProduct);
    assign nxtChkProduct = op1[31:0] * op2[31:0]; 

    always @(posedge clk) begin 
        if ( op2 === 256) begin
            if (~fail)
                $display("SUCESS\n"); 
            $finish; 
        end
        if ( ~(chkProduct === Product) ) begin 
            $display("%d*%d=%d ACTUAL %d",op1,op2,Product,chkProduct);
            $display("FAILURE\n");
            fail <= 1; 
            $finish;
        end
        //$display("%d*%d=%d\n",op1-1,op2,Product);
    end
endmodule 

module multipler (
    input  [31:0]  op0,
    input  [31:0]  op1,
    output [63:0]  res 
);
wire [5:0] P[63:0];
wire [31:0] p0,p1 ,p2 ,p3 ,p4 ,p5 ,p6 ,p7 ,p8 ,p9 ,p10 ,p11 ,p12 ,p13 ,p14 ,p15 ,p16 ,p17 ,p18 ,p19 ,p20 ,p21 ,p22 ,p23 ,p24 ,p25 ,p26 ,p27 ,p28 ,p29 ,p30 ,p31 ;
assign p0[31:0] = {32{op0[0]}} & op1[31:0];
assign p1[31:0] = {32{op0[1]}} & op1[31:0];
assign p2[31:0] = {32{op0[2]}} & op1[31:0];
assign p3[31:0] = {32{op0[3]}} & op1[31:0];
assign p4[31:0] = {32{op0[4]}} & op1[31:0];
assign p5[31:0] = {32{op0[5]}} & op1[31:0];
assign p6[31:0] = {32{op0[6]}} & op1[31:0];
assign p7[31:0] = {32{op0[7]}} & op1[31:0];
assign p8[31:0] = {32{op0[8]}} & op1[31:0];
assign p9[31:0] = {32{op0[9]}} & op1[31:0];
assign p10[31:0] = {32{op0[10]}} & op1[31:0];
assign p11[31:0] = {32{op0[11]}} & op1[31:0];
assign p12[31:0] = {32{op0[12]}} & op1[31:0];
assign p13[31:0] = {32{op0[13]}} & op1[31:0];
assign p14[31:0] = {32{op0[14]}} & op1[31:0];
assign p15[31:0] = {32{op0[15]}} & op1[31:0];
assign p16[31:0] = {32{op0[16]}} & op1[31:0];
assign p17[31:0] = {32{op0[17]}} & op1[31:0];
assign p18[31:0] = {32{op0[18]}} & op1[31:0];
assign p19[31:0] = {32{op0[19]}} & op1[31:0];
assign p20[31:0] = {32{op0[20]}} & op1[31:0];
assign p21[31:0] = {32{op0[21]}} & op1[31:0];
assign p22[31:0] = {32{op0[22]}} & op1[31:0];
assign p23[31:0] = {32{op0[23]}} & op1[31:0];
assign p24[31:0] = {32{op0[24]}} & op1[31:0];
assign p25[31:0] = {32{op0[25]}} & op1[31:0];
assign p26[31:0] = {32{op0[26]}} & op1[31:0];
assign p27[31:0] = {32{op0[27]}} & op1[31:0];
assign p28[31:0] = {32{op0[28]}} & op1[31:0];
assign p29[31:0] = {32{op0[29]}} & op1[31:0];
assign p30[31:0] = {32{op0[30]}} & op1[31:0];
assign p31[31:0] = {32{op0[31]}} & op1[31:0];
assign P[0] = p0[0] +  0;
assign P[1] = p0[1] +  p1[0] + P[0][5:1];
assign P[2] = p0[2] +  p1[1] +  p2[0] + P[1][5:1];
assign P[3] = p0[3] +  p1[2] +  p2[1] +  p3[0] + P[2][5:1];
assign P[4] = p0[4] +  p1[3] +  p2[2] +  p3[1] +  p4[0] + P[3][5:1];
assign P[5] = p0[5] +  p1[4] +  p2[3] +  p3[2] +  p4[1] +  p5[0] + P[4][5:1];
assign P[6] = p0[6] +  p1[5] +  p2[4] +  p3[3] +  p4[2] +  p5[1] +  p6[0] + P[5][5:1];
assign P[7] = p0[7] +  p1[6] +  p2[5] +  p3[4] +  p4[3] +  p5[2] +  p6[1] +  p7[0] + P[6][5:1];
assign P[8] = p0[8] +  p1[7] +  p2[6] +  p3[5] +  p4[4] +  p5[3] +  p6[2] +  p7[1] +  p8[0] + P[7][5:1];
assign P[9] = p0[9] +  p1[8] +  p2[7] +  p3[6] +  p4[5] +  p5[4] +  p6[3] +  p7[2] +  p8[1] +  p9[0] + P[8][5:1];
assign P[10] = p0[10] +  p1[9] +  p2[8] +  p3[7] +  p4[6] +  p5[5] +  p6[4] +  p7[3] +  p8[2] +  p9[1] +  p10[0] + P[9][5:1];
assign P[11] = p0[11] +  p1[10] +  p2[9] +  p3[8] +  p4[7] +  p5[6] +  p6[5] +  p7[4] +  p8[3] +  p9[2] +  p10[1] +  p11[0] + P[10][5:1];
assign P[12] = p0[12] +  p1[11] +  p2[10] +  p3[9] +  p4[8] +  p5[7] +  p6[6] +  p7[5] +  p8[4] +  p9[3] +  p10[2] +  p11[1] +  p12[0] + P[11][5:1];
assign P[13] = p0[13] +  p1[12] +  p2[11] +  p3[10] +  p4[9] +  p5[8] +  p6[7] +  p7[6] +  p8[5] +  p9[4] +  p10[3] +  p11[2] +  p12[1] +  p13[0] + P[12][5:1];
assign P[14] = p0[14] +  p1[13] +  p2[12] +  p3[11] +  p4[10] +  p5[9] +  p6[8] +  p7[7] +  p8[6] +  p9[5] +  p10[4] +  p11[3] +  p12[2] +  p13[1] +  p14[0] + P[13][5:1];
assign P[15] = p0[15] +  p1[14] +  p2[13] +  p3[12] +  p4[11] +  p5[10] +  p6[9] +  p7[8] +  p8[7] +  p9[6] +  p10[5] +  p11[4] +  p12[3] +  p13[2] +  p14[1] +  p15[0] + P[14][5:1];
assign P[16] = p0[16] +  p1[15] +  p2[14] +  p3[13] +  p4[12] +  p5[11] +  p6[10] +  p7[9] +  p8[8] +  p9[7] +  p10[6] +  p11[5] +  p12[4] +  p13[3] +  p14[2] +  p15[1] +  p16[0] + P[15][5:1];
assign P[17] = p0[17] +  p1[16] +  p2[15] +  p3[14] +  p4[13] +  p5[12] +  p6[11] +  p7[10] +  p8[9] +  p9[8] +  p10[7] +  p11[6] +  p12[5] +  p13[4] +  p14[3] +  p15[2] +  p16[1] +  p17[0] + P[16][5:1];
assign P[18] = p0[18] +  p1[17] +  p2[16] +  p3[15] +  p4[14] +  p5[13] +  p6[12] +  p7[11] +  p8[10] +  p9[9] +  p10[8] +  p11[7] +  p12[6] +  p13[5] +  p14[4] +  p15[3] +  p16[2] +  p17[1] +  p18[0] + P[17][5:1];
assign P[19] = p0[19] +  p1[18] +  p2[17] +  p3[16] +  p4[15] +  p5[14] +  p6[13] +  p7[12] +  p8[11] +  p9[10] +  p10[9] +  p11[8] +  p12[7] +  p13[6] +  p14[5] +  p15[4] +  p16[3] +  p17[2] +  p18[1] +  p19[0] + P[18][5:1];
assign P[20] = p0[20] +  p1[19] +  p2[18] +  p3[17] +  p4[16] +  p5[15] +  p6[14] +  p7[13] +  p8[12] +  p9[11] +  p10[10] +  p11[9] +  p12[8] +  p13[7] +  p14[6] +  p15[5] +  p16[4] +  p17[3] +  p18[2] +  p19[1] +  p20[0] + P[19][5:1];
assign P[21] = p0[21] +  p1[20] +  p2[19] +  p3[18] +  p4[17] +  p5[16] +  p6[15] +  p7[14] +  p8[13] +  p9[12] +  p10[11] +  p11[10] +  p12[9] +  p13[8] +  p14[7] +  p15[6] +  p16[5] +  p17[4] +  p18[3] +  p19[2] +  p20[1] +  p21[0] + P[20][5:1];
assign P[22] = p0[22] +  p1[21] +  p2[20] +  p3[19] +  p4[18] +  p5[17] +  p6[16] +  p7[15] +  p8[14] +  p9[13] +  p10[12] +  p11[11] +  p12[10] +  p13[9] +  p14[8] +  p15[7] +  p16[6] +  p17[5] +  p18[4] +  p19[3] +  p20[2] +  p21[1] +  p22[0] + P[21][5:1];
assign P[23] = p0[23] +  p1[22] +  p2[21] +  p3[20] +  p4[19] +  p5[18] +  p6[17] +  p7[16] +  p8[15] +  p9[14] +  p10[13] +  p11[12] +  p12[11] +  p13[10] +  p14[9] +  p15[8] +  p16[7] +  p17[6] +  p18[5] +  p19[4] +  p20[3] +  p21[2] +  p22[1] +  p23[0] + P[22][5:1];
assign P[24] = p0[24] +  p1[23] +  p2[22] +  p3[21] +  p4[20] +  p5[19] +  p6[18] +  p7[17] +  p8[16] +  p9[15] +  p10[14] +  p11[13] +  p12[12] +  p13[11] +  p14[10] +  p15[9] +  p16[8] +  p17[7] +  p18[6] +  p19[5] +  p20[4] +  p21[3] +  p22[2] +  p23[1] +  p24[0] + P[23][5:1];
assign P[25] = p0[25] +  p1[24] +  p2[23] +  p3[22] +  p4[21] +  p5[20] +  p6[19] +  p7[18] +  p8[17] +  p9[16] +  p10[15] +  p11[14] +  p12[13] +  p13[12] +  p14[11] +  p15[10] +  p16[9] +  p17[8] +  p18[7] +  p19[6] +  p20[5] +  p21[4] +  p22[3] +  p23[2] +  p24[1] +  p25[0] + P[24][5:1];
assign P[26] = p0[26] +  p1[25] +  p2[24] +  p3[23] +  p4[22] +  p5[21] +  p6[20] +  p7[19] +  p8[18] +  p9[17] +  p10[16] +  p11[15] +  p12[14] +  p13[13] +  p14[12] +  p15[11] +  p16[10] +  p17[9] +  p18[8] +  p19[7] +  p20[6] +  p21[5] +  p22[4] +  p23[3] +  p24[2] +  p25[1] +  p26[0] + P[25][5:1];
assign P[27] = p0[27] +  p1[26] +  p2[25] +  p3[24] +  p4[23] +  p5[22] +  p6[21] +  p7[20] +  p8[19] +  p9[18] +  p10[17] +  p11[16] +  p12[15] +  p13[14] +  p14[13] +  p15[12] +  p16[11] +  p17[10] +  p18[9] +  p19[8] +  p20[7] +  p21[6] +  p22[5] +  p23[4] +  p24[3] +  p25[2] +  p26[1] +  p27[0] + P[26][5:1];
assign P[28] = p0[28] +  p1[27] +  p2[26] +  p3[25] +  p4[24] +  p5[23] +  p6[22] +  p7[21] +  p8[20] +  p9[19] +  p10[18] +  p11[17] +  p12[16] +  p13[15] +  p14[14] +  p15[13] +  p16[12] +  p17[11] +  p18[10] +  p19[9] +  p20[8] +  p21[7] +  p22[6] +  p23[5] +  p24[4] +  p25[3] +  p26[2] +  p27[1] +  p28[0] + P[27][5:1];
assign P[29] = p0[29] +  p1[28] +  p2[27] +  p3[26] +  p4[25] +  p5[24] +  p6[23] +  p7[22] +  p8[21] +  p9[20] +  p10[19] +  p11[18] +  p12[17] +  p13[16] +  p14[15] +  p15[14] +  p16[13] +  p17[12] +  p18[11] +  p19[10] +  p20[9] +  p21[8] +  p22[7] +  p23[6] +  p24[5] +  p25[4] +  p26[3] +  p27[2] +  p28[1] +  p29[0] + P[28][5:1];
assign P[30] = p0[30] +  p1[29] +  p2[28] +  p3[27] +  p4[26] +  p5[25] +  p6[24] +  p7[23] +  p8[22] +  p9[21] +  p10[20] +  p11[19] +  p12[18] +  p13[17] +  p14[16] +  p15[15] +  p16[14] +  p17[13] +  p18[12] +  p19[11] +  p20[10] +  p21[9] +  p22[8] +  p23[7] +  p24[6] +  p25[5] +  p26[4] +  p27[3] +  p28[2] +  p29[1] +  p30[0] + P[29][5:1];
assign P[31] = p0[31] +  p1[30] +  p2[29] +  p3[28] +  p4[27] +  p5[26] +  p6[25] +  p7[24] +  p8[23] +  p9[22] +  p10[21] +  p11[20] +  p12[19] +  p13[18] +  p14[17] +  p15[16] +  p16[15] +  p17[14] +  p18[13] +  p19[12] +  p20[11] +  p21[10] +  p22[9] +  p23[8] +  p24[7] +  p25[6] +  p26[5] +  p27[4] +  p28[3] +  p29[2] +  p30[1] +  p31[0] + P[30][5:1];
assign P[32] = p1[31] +  p2[30] +  p3[29] +  p4[28] +  p5[27] +  p6[26] +  p7[25] +  p8[24] +  p9[23] +  p10[22] +  p11[21] +  p12[20] +  p13[19] +  p14[18] +  p15[17] +  p16[16] +  p17[15] +  p18[14] +  p19[13] +  p20[12] +  p21[11] +  p22[10] +  p23[9] +  p24[8] +  p25[7] +  p26[6] +  p27[5] +  p28[4] +  p29[3] +  p30[2] +  p31[1] + P[31][5:1];
assign P[33] = p2[31] +  p3[30] +  p4[29] +  p5[28] +  p6[27] +  p7[26] +  p8[25] +  p9[24] +  p10[23] +  p11[22] +  p12[21] +  p13[20] +  p14[19] +  p15[18] +  p16[17] +  p17[16] +  p18[15] +  p19[14] +  p20[13] +  p21[12] +  p22[11] +  p23[10] +  p24[9] +  p25[8] +  p26[7] +  p27[6] +  p28[5] +  p29[4] +  p30[3] +  p31[2] + P[32][5:1];
assign P[34] = p3[31] +  p4[30] +  p5[29] +  p6[28] +  p7[27] +  p8[26] +  p9[25] +  p10[24] +  p11[23] +  p12[22] +  p13[21] +  p14[20] +  p15[19] +  p16[18] +  p17[17] +  p18[16] +  p19[15] +  p20[14] +  p21[13] +  p22[12] +  p23[11] +  p24[10] +  p25[9] +  p26[8] +  p27[7] +  p28[6] +  p29[5] +  p30[4] +  p31[3] + P[33][5:1];
assign P[35] = p4[31] +  p5[30] +  p6[29] +  p7[28] +  p8[27] +  p9[26] +  p10[25] +  p11[24] +  p12[23] +  p13[22] +  p14[21] +  p15[20] +  p16[19] +  p17[18] +  p18[17] +  p19[16] +  p20[15] +  p21[14] +  p22[13] +  p23[12] +  p24[11] +  p25[10] +  p26[9] +  p27[8] +  p28[7] +  p29[6] +  p30[5] +  p31[4] + P[34][5:1];
assign P[36] = p5[31] +  p6[30] +  p7[29] +  p8[28] +  p9[27] +  p10[26] +  p11[25] +  p12[24] +  p13[23] +  p14[22] +  p15[21] +  p16[20] +  p17[19] +  p18[18] +  p19[17] +  p20[16] +  p21[15] +  p22[14] +  p23[13] +  p24[12] +  p25[11] +  p26[10] +  p27[9] +  p28[8] +  p29[7] +  p30[6] +  p31[5] + P[35][5:1];
assign P[37] = p6[31] +  p7[30] +  p8[29] +  p9[28] +  p10[27] +  p11[26] +  p12[25] +  p13[24] +  p14[23] +  p15[22] +  p16[21] +  p17[20] +  p18[19] +  p19[18] +  p20[17] +  p21[16] +  p22[15] +  p23[14] +  p24[13] +  p25[12] +  p26[11] +  p27[10] +  p28[9] +  p29[8] +  p30[7] +  p31[6] + P[36][5:1];
assign P[38] = p7[31] +  p8[30] +  p9[29] +  p10[28] +  p11[27] +  p12[26] +  p13[25] +  p14[24] +  p15[23] +  p16[22] +  p17[21] +  p18[20] +  p19[19] +  p20[18] +  p21[17] +  p22[16] +  p23[15] +  p24[14] +  p25[13] +  p26[12] +  p27[11] +  p28[10] +  p29[9] +  p30[8] +  p31[7] + P[37][5:1];
assign P[39] = p8[31] +  p9[30] +  p10[29] +  p11[28] +  p12[27] +  p13[26] +  p14[25] +  p15[24] +  p16[23] +  p17[22] +  p18[21] +  p19[20] +  p20[19] +  p21[18] +  p22[17] +  p23[16] +  p24[15] +  p25[14] +  p26[13] +  p27[12] +  p28[11] +  p29[10] +  p30[9] +  p31[8] + P[38][5:1];
assign P[40] = p9[31] +  p10[30] +  p11[29] +  p12[28] +  p13[27] +  p14[26] +  p15[25] +  p16[24] +  p17[23] +  p18[22] +  p19[21] +  p20[20] +  p21[19] +  p22[18] +  p23[17] +  p24[16] +  p25[15] +  p26[14] +  p27[13] +  p28[12] +  p29[11] +  p30[10] +  p31[9] + P[39][5:1];
assign P[41] = p10[31] +  p11[30] +  p12[29] +  p13[28] +  p14[27] +  p15[26] +  p16[25] +  p17[24] +  p18[23] +  p19[22] +  p20[21] +  p21[20] +  p22[19] +  p23[18] +  p24[17] +  p25[16] +  p26[15] +  p27[14] +  p28[13] +  p29[12] +  p30[11] +  p31[10] + P[40][5:1];
assign P[42] = p11[31] +  p12[30] +  p13[29] +  p14[28] +  p15[27] +  p16[26] +  p17[25] +  p18[24] +  p19[23] +  p20[22] +  p21[21] +  p22[20] +  p23[19] +  p24[18] +  p25[17] +  p26[16] +  p27[15] +  p28[14] +  p29[13] +  p30[12] +  p31[11] + P[41][5:1];
assign P[43] = p12[31] +  p13[30] +  p14[29] +  p15[28] +  p16[27] +  p17[26] +  p18[25] +  p19[24] +  p20[23] +  p21[22] +  p22[21] +  p23[20] +  p24[19] +  p25[18] +  p26[17] +  p27[16] +  p28[15] +  p29[14] +  p30[13] +  p31[12] + P[42][5:1];
assign P[44] = p13[31] +  p14[30] +  p15[29] +  p16[28] +  p17[27] +  p18[26] +  p19[25] +  p20[24] +  p21[23] +  p22[22] +  p23[21] +  p24[20] +  p25[19] +  p26[18] +  p27[17] +  p28[16] +  p29[15] +  p30[14] +  p31[13] + P[43][5:1];
assign P[45] = p14[31] +  p15[30] +  p16[29] +  p17[28] +  p18[27] +  p19[26] +  p20[25] +  p21[24] +  p22[23] +  p23[22] +  p24[21] +  p25[20] +  p26[19] +  p27[18] +  p28[17] +  p29[16] +  p30[15] +  p31[14] + P[44][5:1];
assign P[46] = p15[31] +  p16[30] +  p17[29] +  p18[28] +  p19[27] +  p20[26] +  p21[25] +  p22[24] +  p23[23] +  p24[22] +  p25[21] +  p26[20] +  p27[19] +  p28[18] +  p29[17] +  p30[16] +  p31[15] + P[45][5:1];
assign P[47] = p16[31] +  p17[30] +  p18[29] +  p19[28] +  p20[27] +  p21[26] +  p22[25] +  p23[24] +  p24[23] +  p25[22] +  p26[21] +  p27[20] +  p28[19] +  p29[18] +  p30[17] +  p31[16] + P[46][5:1];
assign P[48] = p17[31] +  p18[30] +  p19[29] +  p20[28] +  p21[27] +  p22[26] +  p23[25] +  p24[24] +  p25[23] +  p26[22] +  p27[21] +  p28[20] +  p29[19] +  p30[18] +  p31[17] + P[47][5:1];
assign P[49] = p18[31] +  p19[30] +  p20[29] +  p21[28] +  p22[27] +  p23[26] +  p24[25] +  p25[24] +  p26[23] +  p27[22] +  p28[21] +  p29[20] +  p30[19] +  p31[18] + P[48][5:1];
assign P[50] = p19[31] +  p20[30] +  p21[29] +  p22[28] +  p23[27] +  p24[26] +  p25[25] +  p26[24] +  p27[23] +  p28[22] +  p29[21] +  p30[20] +  p31[19] + P[49][5:1];
assign P[51] = p20[31] +  p21[30] +  p22[29] +  p23[28] +  p24[27] +  p25[26] +  p26[25] +  p27[24] +  p28[23] +  p29[22] +  p30[21] +  p31[20] + P[50][5:1];
assign P[52] = p21[31] +  p22[30] +  p23[29] +  p24[28] +  p25[27] +  p26[26] +  p27[25] +  p28[24] +  p29[23] +  p30[22] +  p31[21] + P[51][5:1];
assign P[53] = p22[31] +  p23[30] +  p24[29] +  p25[28] +  p26[27] +  p27[26] +  p28[25] +  p29[24] +  p30[23] +  p31[22] + P[52][5:1];
assign P[54] = p23[31] +  p24[30] +  p25[29] +  p26[28] +  p27[27] +  p28[26] +  p29[25] +  p30[24] +  p31[23] + P[53][5:1];
assign P[55] = p24[31] +  p25[30] +  p26[29] +  p27[28] +  p28[27] +  p29[26] +  p30[25] +  p31[24] + P[54][5:1];
assign P[56] = p25[31] +  p26[30] +  p27[29] +  p28[28] +  p29[27] +  p30[26] +  p31[25] + P[55][5:1];
assign P[57] = p26[31] +  p27[30] +  p28[29] +  p29[28] +  p30[27] +  p31[26] + P[56][5:1];
assign P[58] = p27[31] +  p28[30] +  p29[29] +  p30[28] +  p31[27] + P[57][5:1];
assign P[59] = p28[31] +  p29[30] +  p30[29] +  p31[28] + P[58][5:1];
assign P[60] = p29[31] +  p30[30] +  p31[29] + P[59][5:1];
assign P[61] = p30[31] +  p31[30] + P[60][5:1];
assign P[62] = p31[31] + P[61][5:1];
assign P[63] =P[62][5:1];
assign       res[63:0] = {P[63][0],P[62][0],P[61][0],P[60][0],P[59][0],P[58][0],P[57][0],P[56][0],P[55][0],P[54][0],P[53][0],P[52][0],P[51][0],P[50][0],P[49][0],P[48][0],P[47][0],P[46][0],P[45][0],P[44][0],P[43][0],P[42][0],P[41][0],P[40][0],P[39][0],P[38][0],P[37][0],P[36][0],P[35][0],P[34][0],P[33][0],P[32][0],P[31][0],P[30][0],P[29][0],P[28][0],P[27][0],P[26][0],P[25][0],P[24][0],P[23][0],P[22][0],P[21][0],P[20][0],P[19][0],P[18][0],P[17][0],P[16][0],P[15][0],P[14][0],P[13][0],P[12][0],P[11][0],P[10][0],P[9][0],P[8][0],P[7][0],P[6][0],P[5][0],P[4][0],P[3][0],P[2][0],P[1][0],P[0][0]};
endmodule
